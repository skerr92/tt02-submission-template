module shiftreg
  ( input wire decode[3:0],
   input wire clk, reset, data_in,
   output wire data_out[7:0]
  );
  
  always @(posedge clk) begin
    
  end
endmodule
